
//iverilog -o "helloworld.vvp" helloworld.v
//vvp helloworld.vvp

module helloworld ;

initial begin
    $display("hello , world!");
end
    
endmodule